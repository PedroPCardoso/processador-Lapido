module banco_registrador_tb();





endmodule
