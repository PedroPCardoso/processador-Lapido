library verilog;
use verilog.vl_types.all;
entity registerFile_tb is
end registerFile_tb;
