// inicializa o dispositivo e passa o controle para a Unidade de Controle
module bios (CLK);
input CLK;
input [31:0] D;
output [31:0] Q;
reg [31:0] Q;

	always @(posedge CLK)
	begin
		// Carrega memória
		// Inicializa valores dos componentes
	end
			
endmodule