module ULA_TB();

  reg [31:0] a, b;
  wire flag;
  wire [31:0] out;
  reg [4:0] opcode;


   ULA ULA(
      .A(a),
      .B(b),
      .opcode(opcode),
      .Flag(flag),
      .Out(out)
      );

    initial begin
      a=32'b00000000000000000000000000000001;
      b=32'b00000000000000000000000000000000;
      opcode=5'b0000;
      $display(out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000011;
      opcode=5'b00001;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000011;
      opcode=5'b00011;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000011;
      opcode=5'b00100;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000011;
      opcode=5'b00101;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000011;
      opcode=5'b00110;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b01000;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b01001;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b10000;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b10001;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b10010;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b10011;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b10100;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b10101;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b10110;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b10111;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b11000;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b11001;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b11010;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b11011;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b11100;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b11101;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b11110;
      $display (out);

      #100 ;
      a=32'b00000000000000000000000000000101;
      b=32'b00000000000000000000000000000000;
      opcode=5'b11111;
      $display (out);

      end

endmodule
