library verilog;
use verilog.vl_types.all;
entity clockFSM is
end clockFSM;
