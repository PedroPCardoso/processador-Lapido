library verilog;
use verilog.vl_types.all;
entity ULA_TB is
end ULA_TB;
